`define MODULE_NAME Customized_PHY_Top
`define Q0_LN0
`define Q0_LN0_PMA_WIDTH 10
`define Q0_LN0_TX_GEARBOX 1
`define Q0_LN0_RX_GEARBOX 1
`define Q0_LN0_8B10B_ENCODE
`define Q0_LN0_CHANNEL_BONDING_MASTER_SEL 0
`define Q0_LN0_TX_IF_MST_SEL 0
